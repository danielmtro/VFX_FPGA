module inversion_filter_tb;

endmodule 