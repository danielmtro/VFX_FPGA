// scaling.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module scaling (
		input  wire        clk_clk,             //   clk.clk
		input  wire        reset_reset,         // reset.reset
		input  wire        sauce_ready,         // sauce.ready
		output wire        sauce_startofpacket, //      .startofpacket
		output wire        sauce_endofpacket,   //      .endofpacket
		output wire        sauce_valid,         //      .valid
		output wire [11:0] sauce_data,          //      .data
		output wire [1:0]  sauce_channel,       //      .channel
		input  wire        sink_startofpacket,  //  sink.startofpacket
		input  wire        sink_endofpacket,    //      .endofpacket
		input  wire        sink_valid,          //      .valid
		output wire        sink_ready,          //      .ready
		input  wire [11:0] sink_data            //      .data
	);

	scaling_video_scaler_0 video_scaler_0 (
		.clk                      (clk_clk),             //                  clk.clk
		.reset                    (reset_reset),         //                reset.reset
		.stream_in_startofpacket  (sink_startofpacket),  //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (sink_endofpacket),    //                     .endofpacket
		.stream_in_valid          (sink_valid),          //                     .valid
		.stream_in_ready          (sink_ready),          //                     .ready
		.stream_in_data           (sink_data),           //                     .data
		.stream_out_ready         (sauce_ready),         // avalon_scaler_source.ready
		.stream_out_startofpacket (sauce_startofpacket), //                     .startofpacket
		.stream_out_endofpacket   (sauce_endofpacket),   //                     .endofpacket
		.stream_out_valid         (sauce_valid),         //                     .valid
		.stream_out_data          (sauce_data),          //                     .data
		.stream_out_channel       (sauce_channel)        //                     .channel
	);

endmodule
