module data_expander_tb;

endmodule 