//module filter_select_tb;
//
//
//
//
//
//	filter_select DUT(
//	.clk,
//	.reset,
//	.freq_flag,
//	.filter_num,
//	
//
//	.data_in,
//	.sop_in,
//	.eop_in,
//	.valid_in,
//	
//
//	.ready_in,
//
//	.ready_out,
//
//	.data_out,
//	.sop_out,
//	.eop_out,
//	.valid_out) 
//
//
//
//
//
//endmodule 