
module vga_clock (
	clk_clk,
	reset_reset_n,
	vga_clk_clk,
	reset_source_reset);	

	input		clk_clk;
	input		reset_reset_n;
	output		vga_clk_clk;
	output		reset_source_reset;
endmodule
