module filter_select_tb;


endmodule 